`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.02.2025 09:29:41
// Design Name: 
// Module Name: exp4_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module exp4_tb( );
    logic [1:0] a;
    logic [1:0] b;
    logic R, G, B;
exp4 zain (
    .a(a),
    .b(b),
    .R(R),
    .G(G),
    .B(B)
);
initial begin
        a[1]=0; a[0]=0; b[1]=0 ; b[0]=0;
        #10;
        a[1]=0; a[0]=0; b[1]=0 ; b[0]=1;
        #10;
        a[1]=0; a[0]=0; b[1]=1 ; b[0]=0;
        #10;
        a[1]=0; a[0]=0; b[1]=1 ; b[0]=1;
        #10;
        a[1]=0; a[0]=1; b[1]=0 ; b[0]=0;
        #10;
        a[1]=0; a[0]=1; b[1]=0 ; b[0]=1;
        #10;
        a[1]=0; a[0]=1; b[1]=1 ; b[0]=0;
        #10;
        a[1]=0; a[0]=1; b[1]=1 ; b[0]=1;
        #10;
        a[1]=1; a[0]=0; b[1]=0 ; b[0]=0;
        #10;
        a[1]=1; a[0]=0; b[1]=0 ; b[0]=1;
        #10;
        a[1]=1; a[0]=0; b[1]=1 ; b[0]=0;
        #10;
        a[1]=1; a[0]=0; b[1]=1 ; b[0]=1;
        #10;
        a[1]=1; a[0]=1; b[1]=0 ; b[0]=0;
        #10;
        a[1]=1; a[0]=1; b[1]=0 ; b[0]=1;
        #10;
        a[1]=1; a[0]=1; b[1]=1 ; b[0]=0;
        #10;
        a[1]=1; a[0]=1; b[1]=1 ; b[0]=1;
        #10;
        $stop;
        end    

    
endmodule
